module valid_result(
    input wire valid_address,
    output wire valid_result
);
    assign valid_result = valid_address;
endmodule